/*
Guia_0103a - Arquitetura de computadores
Autor: Izadora Galarza Alves
*/

module guia_0103d;

integer x=157;
reg[7:0] b=0;

initial
begin:main

$display("Guia_0103 - D");
$display("X= %d",x);
$display("b=%8b",b);
b=x;
$display("b= %8b(2) / %o(8) / %x(16)",b,b,b);

end
endmodule